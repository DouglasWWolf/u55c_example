//================================================================================================
//    Date      Vers   Who  Changes
// -----------------------------------------------------------------------------------------------
// 04-Jun-2025  1.0.0  DWW  Initial creation
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;
localparam RTL_TYPE      = 60425;
localparam RTL_SUBTYPE   = 0;

localparam VERSION_DAY   = 4;
localparam VERSION_MONTH = 6;
localparam VERSION_YEAR  = 2025;
